module Test_bench_of_Signed_Calculator_4bit();

reg A3, A2, A1, A0, B3, B2, B1, B0, M1, M0, S1, S0, Reset;
wire Out15_R7, Out14_R6, Out13_R5, Out12_R4, Out11_R3, Out10_R2, Out9_R1, Out8_R0, Out7, Out6, Out5, Out4, Out3, Out2, Out1, Out0;

Signed_Calculator_4bit_Reset DUT(Out15_R7, Out14_R6, Out13_R5, Out12_R4, Out11_R3, Out10_R2, Out9_R1, Out8_R0, Out7, Out6, Out5, Out4, Out3, Out2, Out1, Out0, A3, A2, A1, A0, B3, B2, B1, B0, M1, M0, S1, S0, Reset);

initial
begin

Reset =1'b0; A3= 1'b1; A2= 1'b0; A1=1'b1; A0=1'b0; B3= 1'b0; B2= 1'b1; B1= 1'b1; B0=1'b1; M1= 1'b0; M0= 1'b1; S1= 1'b1; S0= 1'b1;
#1 M1= 1'b1; M0= 1'b1; 
#1 A3= 1'b0; A1= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0; 

Reset = 1'b1;
M1= 1'b0; M0= 1'b0;  // Addition of +A +B

#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

//////////////////////Addition of +A -B ////////////////////

S1= 1'b1; S0= 1'b0;

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

/////////////////////////Addition of -A +B /////////////////////////////////////

#1 S1= 1'b0; S0= 1'b1; 

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

/////////////////////////Addition of -A -B /////////////////////////////////////

#1 S1= 1'b0; S0= 1'b0; 

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

///////////////////////////////////Subtraction of +A +B////////////////////////////////////

M1= 1'b0; M0= 1'b1;


#1 S1=1'b1; S0= 1'b1;

A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

//////////////////////Subtraction of +A -B ////////////////////

S1= 1'b1; S0= 1'b0;

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

/////////////////////////Subtraction of -A +B /////////////////////////////////////

#1 S1= 1'b0; S0= 1'b1; 

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

/////////////////////////Subtraction of -A -B /////////////////////////////////////

#1 S1= 1'b0; S0= 1'b0; 

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 


///////////////////////////////////Multiplication of +A +B////////////////////////////////////

M1= 1'b1; M0= 1'b0;


#1 S1=1'b1; S0= 1'b1;

A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

//////////////////////Multiplication of +A -B ////////////////////

S1= 1'b1; S0= 1'b0;

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

/////////////////////////Multiplication of -A +B /////////////////////////////////////

#1 S1= 1'b0; S0= 1'b1; 

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

/////////////////////////Multiplication of -A -B /////////////////////////////////////

#1 S1= 1'b0; S0= 1'b0; 

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 


///////////////////////////////////Division of +A +B////////////////////////////////////

M1= 1'b1; M0= 1'b1;


#1 S1=1'b1; S0= 1'b1;

A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

//////////////////////Division of +A -B ////////////////////

S1= 1'b1; S0= 1'b0;

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

/////////////////////////Division of -A +B /////////////////////////////////////

#1 S1= 1'b0; S0= 1'b1; 

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

/////////////////////////Division of -A -B /////////////////////////////////////

#1 S1= 1'b0; S0= 1'b0; 

#1 A3= 1'b0; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3= 1'b0; B2= 1'b0; B1= 1'b0; B0= 1'b0;
#1 B0=1'b1;  // A=0, B= 0-->15 
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=1, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=2, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=3, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=4, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=5, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=6, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=7, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A3= 1'b1; A2= 1'b0; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=8, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=9, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=10, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b0; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=11, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=12, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b0; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=13, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b0; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=14, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 

#1 A2= 1'b1; A1= 1'b1; A0= 1'b1; B3=1'b0; B2=1'b0; B1=1'b0; B0=1'b0; // A=15, B= 0-->15
#1 B0=1'b1;   
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B3=1'b1; B2=1'b0; B1=1'b0; B0=1'b0;
#1 B0=1'b1;  
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1;
#1 B2= 1'b1; B1=1'b0; B0=1'b0;
#1 B0=1'b1;
#1 B1=1'b1; B0=1'b0;
#1 B0=1'b1; 



#1 $finish;
end
endmodule
